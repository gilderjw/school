// Verilog test fixture created from schematic /home/wangs4/1516a-csse232-sid-transputer/XilinxProject/ALU-praise be unto him/Test_ALUMem.sch - Tue Nov  3 18:48:49 2015

`timescale 1ns / 1ps

module Test_ALUMem_Test_ALUMem_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Test_ALUMem UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
